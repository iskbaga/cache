module address();

reg [9:0] tag [0:7807];
reg [9:0] index [0:7807];
reg [9:0] offset [0:7807]; 

endmodule