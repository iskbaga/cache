module ram();

parameter size = 4096; 

reg [127:0] ram [0:size-1]; 

endmodule